-- Laboratory RA solutions/versuch1
-- Sommersemester 24
-- Group Details
-- Lab Date:
-- 1. Participant First and Last Name: 
-- 2. Participant First and Last Name:


library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;
  use ieee.math_real.all;
  use work.constant_package.all;

entity gen_mux_tb is
end entity gen_mux_tb;

architecture behavior of gen_mux_tb is
-- begin solution:
 -- end solution!!
end architecture behavior;