-- Laboratory RA solutions/versuch2
-- Sommersemester 24
-- Group Details
-- Lab Date:
-- 1. Participant First and Last Name: 
-- 2. Participant First and Last Name:

library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;
  use ieee.math_real.all;
  use work.constant_package.all;

entity register_file is
-- begin solution:
   -- end solution!!
end entity register_file;

architecture arc of register_file is
-- begin solution:
   -- end solution!!
end architecture arc;
