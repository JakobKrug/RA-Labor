-- Laboratory RA solutions/versuch1
-- Sommersemester 24
-- Group Details
-- Lab Date:
-- 1. Participant First and Last Name: 
-- 2. Participant First and Last Name:


library ieee;
  use ieee.std_logic_1164.all;
  use work.constant_package.all;

entity gen_mux is
  -- begin solution:
  -- end solution!!
end entity gen_mux;

architecture dataflow of gen_mux is
-- begin solution:
-- end solution!!
end architecture dataflow;
