-- Laboratory RA solutions/versuch1
-- Sommersemester 24
-- Group Details
-- Lab Date:
-- 1. Participant First and Last Name: 
-- 2. Participant First and Last Name:


library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.Constant_Package.all;

entity gen_register_tb is
end entity gen_register_tb;

architecture testbench of gen_register_tb is
-- begin solution:
-- end solution!!
end architecture testbench;